library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.parameter_pkg.all;
use work.types_pkg.all;

entity mem_control is
	generic(
		mem_type : memory_type := P_MEM
	);
	port(
		clk, rst        : in std_logic;
		rd_addr         : in unsigned(BW_ADDRESS-1 downto 0);
		rd_en           : in std_logic;
		data_out        : out std_logic_vector(23 downto 0);
		data_out_valid  : out std_logic;
		wr_addr         : in  unsigned(BW_ADDRESS-1 downto 0);
		wr_en           : in  std_logic;
		wr_accomplished : out std_logic;
		data_in         : in  std_logic_vector(23 downto 0)
	);
end entity mem_control;


architecture rtl of mem_control is

	signal int_mem_rd_addr : std_logic_vector(7 downto 0);
	type int_mem_type is array(0 to 255) of std_logic_vector(23 downto 0);
	signal int_mem : int_mem_type;
	signal int_pmem : int_mem_type := (
-- ABS begin
--X"0000B9",
--X"56F400",
--X"200000",
--X"200026",
--X"56F400",
--X"E00000",
--X"200026",
--X"56F400",
--X"000000",
--X"200026",
--X"52F400",
--X"000080",
--X"200026",
-- ABS end

-- ADC begin
--X"46F400",
--X"000000",
--X"47F400",
--X"000001",
--X"20001B",
--X"51F400",
--X"000001",
--X"0000B9",
--X"0001F9",
--X"200039",
--X"47F400",
--X"800000",
--X"53F400",
--X"000080",
--X"200039",
-- ADC end

-- ADD begin
--X"46F400",
--X"000000",
--X"47F400",
--X"000001",
--X"20001B",
--X"51F400",
--X"000001",
--X"0000B9",
--X"0001F9",
--X"200038",
--X"47F400",
--X"800000",
--X"53F400",
--X"000080",
--X"200038",
-- ADD end

-- ADDL begin
--X"56F400",
--X"000055",
--X"20001B",
--X"51F400",
--X"000055",
--X"0000B9",
--X"20001A",
--X"56F400",
--X"0000AA",
--X"20001A",
--X"53F400",
--X"000080",
--X"20001A",
-- ADDL end

-- ADDR begin
--X"56F400",
--X"000055",
--X"20001B",
--X"51F400",
--X"000055",
--X"0000B9",
--X"20000A",
--X"56F400",
--X"0000AA",
--X"20000A",
--X"53F400",
--X"000080",
--X"20000A",
-- ADDR end

-- AND begin
--X"46F400",
--X"000FFF",
--X"57F400",
--X"FFFFFF",
--X"0000B9",
--X"20005E",
--X"46F400",
--X"FFF000",
--X"57F400",
--X"FFFFFF",
--X"0000B9",
--X"20005E",
--X"46F400",
--X"000000",
--X"57F400",
--X"FFFFFF",
--X"0000B9",
--X"20005E",
-- AND end

-- EOR begin
--X"46F400",
--X"000FFF",
--X"57F400",
--X"FF00FF",
--X"0000B9",
--X"20005B",
--X"46F400",
--X"FFFFFF",
--X"57F400",
--X"FFFFFF",
--X"0000B9",
--X"20005B",
-- EOR end

-- OR begin
--X"46F400",
--X"000FFF",
--X"57F400",
--X"FF00FF",
--X"0000B9",
--X"20005A",
--X"46F400",
--X"000000",
--X"57F400",
--X"000000",
--X"0000B9",
--X"20005A",
-- OR end

-- NOT begin
--X"46F400",
--X"000FFF",
--X"57F400",
--X"7F00FF",
--X"0000B9",
--X"20001F",
--X"46F400",
--X"000000",
--X"57F400",
--X"FFFFFF",
--X"0000B9",
--X"20001F",
-- NOT end

-- ASL begin
--X"20001B",
--X"51F400",
--X"0000A5",
--X"55F400",
--X"0000A5",
--X"53F400",
--X"0000A5",
--X"0000B9",
--X"20003A",
-- ASL end

-- ASR begin
--X"20001B",
--X"51F400",
--X"0000A5",
--X"55F400",
--X"0000A5",
--X"53F400",
--X"0000A5",
--X"0000B9",
--X"20002A",
-- ASR end

-- CLR begin
--X"0000B9",
--X"56F400",
--X"200000",
--X"200013",
--X"56F400",
--X"E00000",
--X"0000B9",
--X"0001F9",
--X"200013",
-- CLR end

-- CMP begin
--X"2F2000",
--X"262400",
--X"0000B9",
--X"20005D",
--X"2F2000",
--X"262000",
--X"0000B9",
--X"20005D",
--X"2F2400",
--X"262000",
--X"0000B9",
--X"20005D",
--X"57F400",
--X"800AAA",
--X"262000",
--X"0000B9",
--X"20005D",
--X"46F400",
--X"800AAA",
--X"2F2000",
--X"0000B9",
--X"20005D",
-- CMP end

-- CMPM begin
--X"2F2000",
--X"262400",
--X"0000B9",
--X"20005F",
--X"2F2000",
--X"262000",
--X"0000B9",
--X"20005F",
--X"2F2400",
--X"262000",
--X"0000B9",
--X"20005F",
--X"57F400",
--X"800AAA",
--X"262000",
--X"0000B9",
--X"20005F",
--X"46F400",
--X"800AAA",
--X"2F2000",
--X"0000B9",
--X"20005F",
-- CMPM end

-- DIV begin
--X"00FEB9",
--X"44F400",
--X"600000",
--X"56F400",
--X"200000",
--X"0618A0",
--X"018040",
--X"210E00",
-- DIV end

-- LSL begin
--X"0000B9",
--X"56F400",
--X"200000",
--X"56F400",
--X"AAAAAA",
--X"50F400",
--X"BCDEFA",
--X"0618A0",
--X"200033",
-- LSL end

-- LSR begin
--X"0000B9",
--X"56F400",
--X"200000",
--X"56F400",
--X"AAAAAA",
--X"50F400",
--X"BCDEFA",
--X"0618A0",
--X"200023",
-- LSR end

-- MPY begin
--X"0000B9",
--X"44F400",
--X"200000",
--X"46F400",
--X"400000",
--X"2000D0",
--X"44F400",
--X"E00000",
--X"46F400",
--X"B9999A",
--X"2000D0",
--X"44F400",
--X"E66666",
--X"46F400",
--X"466666",
--X"2000D0",
--X"44F400",
--X"E66666",
--X"46F400",
--X"466666",
--X"2000D4",
-- MPY end

-- MAC begin
--X"0000B9",
--X"200013",
--X"2A8000",
--X"44F400",
--X"200000",
--X"46F400",
--X"400000",
--X"2000D6",
--X"44F400",
--X"E00000",
--X"46F400",
--X"B9999A",
--X"2000D2",
--X"44F400",
--X"E66666",
--X"46F400",
--X"466666",
--X"2000D2",
--X"44F400",
--X"E66666",
--X"46F400",
--X"466666",
--X"2000D6",
-- MAC end

-- MACR begin
--X"0000B9",
--X"200013",
--X"2E1000",
--X"44F400",
--X"123456",
--X"46F400",
--X"123456",
--X"2000D3",
--X"56F400",
--X"100001",
--X"44F400",
--X"123456",
--X"46F400",
--X"123456",
--X"2000D3",
--X"2E1000",
--X"50F400",
--X"800000",
--X"44F400",
--X"123456",
--X"46F400",
--X"123456",
--X"2000D3",
-- MACR end

-- MPYR begin
--X"0000B9",
--X"46F400",
--X"654321",
--X"200095",
-- MPYR end

-- NEG begin
--X"0000B9",
--X"56F400",
--X"654321",
--X"200036",
--X"200013",
--X"52F400",
--X"000080",
--X"200036",
--X"56F400",
--X"800000",
--X"200036",
-- NEG end

-- NORM begin
X"200013",
X"2C0100",
X"200003",
X"062FA0",
X"01DB15",
X"200013",
X"2EFF00",
X"2A8400",
X"200003",
X"062FA0",
X"01D915",
X"200013",
X"062FA0",
X"01DA15",
-- NORM end

-- RND begin
--X"0000B9",
--X"54F400",
--X"123456",
--X"50F400",
--X"789ABC",
--X"200011",
--X"54F400",
--X"123456",
--X"50F400",
--X"800000",
--X"200011",
--X"54F400",
--X"123455",
--X"50F400",
--X"800000",
--X"200011",
-- RND end

-- ROR begin
--X"0000B9",
--X"56F400",
--X"AAAAAA",
--X"50F400",
--X"BCDEFA",
--X"0618A0",
--X"200027",
-- ROR end

-- ROL begin
--X"0000B9",
--X"56F400",
--X"AAAAAA",
--X"50F400",
--X"BCDEFA",
--X"0618A0",
--X"200037",
-- ROL end


-- SUB begin
--X"46F400",
--X"000000",
--X"47F400",
--X"000001",
--X"20001B",
--X"51F400",
--X"000001",
--X"0000B9",
--X"0001F9",
--X"20003C",
--X"47F400",
--X"800000",
--X"53F400",
--X"000080",
--X"20003C",
--X"20001B",
--X"53F400",
--X"000080",
--X"47F400",
--X"000001",
--X"20007C",
-- SUB end

-- SUBL begin
--X"50F400",
--X"000000",
--X"54F400",
--X"000001",
--X"20001B",
--X"51F400",
--X"000001",
--X"0000B9",
--X"0001F9",
--X"20001E",
--X"54F400",
--X"800000",
--X"53F400",
--X"000080",
--X"20001E",
--X"20001B",
--X"53F400",
--X"000080",
--X"54F400",
--X"000001",
--X"20001E",
-- SUBL end

-- SUBR begin
--X"50F400",
--X"000000",
--X"54F400",
--X"000001",
--X"20001B",
--X"51F400",
--X"000001",
--X"0000B9",
--X"0001F9",
--X"20000E",
--X"54F400",
--X"800000",
--X"53F400",
--X"000080",
--X"20000E",
--X"20001B",
--X"53F400",
--X"000080",
--X"54F400",
--X"000001",
--X"20000E",
-- SUBR end

-- SBC begin
--X"46F400",
--X"000000",
--X"47F400",
--X"000001",
--X"20001B",
--X"51F400",
--X"000001",
--X"0000B9",
--X"0001F9",
--X"20003D",
--X"47F400",
--X"800000",
--X"53F400",
--X"000080",
--X"20003D",
--X"20001B",
--X"53F400",
--X"000080",
--X"47F400",
--X"000001",
--X"20003D",
-- SBC end

-- TCC begin
--X"311400",
--X"44F400",
--X"ABCDEF",
--X"57F400",
--X"123456",
--X"0000B9",
--X"038143",
--X"03014A",
--X"0004F9",
--X"03A143",
--X"03214A",
-- TCC end

-- TFR begin
--X"56F400",
--X"ABCDEF",
--X"57F400",
--X"123456",
--X"21EE09",
--X"44F400",
--X"555555",
--X"47F400",
--X"AAAAAA",
--X"21C441",
--X"21E679",
-- TFR end

-- TST begin
--X"20001B",
--X"20000B",
--X"0000B9",
--X"0001F9",
--X"53F400",
--X"000080",
--X"20000B",
--X"53F400",
--X"00007F",
--X"20000B",
-- TST end


--X"2AFF00",
--X"54F400",
--X"FFFFFF",
--X"50F400",
--X"FFFFF2",
--X"200026",
--X"000000",
--X"000000",
--X"000000",
--X"000000",
--X"000000",
--X"000000",
--X"000000",
--X"000000",
--X"000000",
--X"000000",
X"000000",
X"000000",
X"000000",
X"000000",
X"000000",
X"000000",
X"000000",
X"000000",
X"000000",
--X"44F400",
--X"100010",
--X"45F400",
--X"100011",
--X"0B5880",
--X"000017",
--X"46F400",
--X"100026",
--X"47F400",
--X"100027",
--X"425800",
--X"435800",
--X"420A00",
--X"431F00",
--X"437000",
--X"0000A0",
--X"427000",
--X"00004F",
--  X"42F800",
--  X"43F800",
--  X"428A00",
--  X"439F00",
--	"001100000100100000000000",  -- 0 move #72,r0
--	"001110000000100000000000",  -- 1 move #8,n0
--	"000001010000000010100000",  -- 2 move #0,m0
--	"000001010001000010100001",  -- 3 move #16,m1
--	"000001101110000100100000",  -- 4 rep m1
--	"010001001100100000000000",  -- 5 move x:(r0)+n0,x0
--	"000000000000000000000000",  -- 6
--	"000000000000000000000000",  -- 7
--	"000000000000000000000000",  -- 8
--	"000000000000000000000000",  -- 9 
--	"000000000000000000000000",  -- 10
--	"000000000000000000000000",  -- 11
--	"000000000000000000000000",  -- 12
--	"000000000000000000000000",  -- 13
--	"000000000000000000000000",  -- 14
--	"000000000000000000000000",  -- 15
--	"000000000000000000000000",  -- 16
--	"000000000000000000000000",  -- 17
--	"000000000000000000000000",  -- 18
--	"000000000000000000000000",  -- 19
--	"000010101101101010000000",  -- 20 -- JMP (r2)+
--	"000000000000000000000000",  -- 20
--	"000000000000000000000000",  -- 21
--	"000000000000000000000000",  -- 22
	"000000000000000000000000",  -- 23
	"000000000000000000000000",  -- 24
	"000000000000000000000000",  -- 25
	"000000000000000000000000",  -- 26
	"000000000000000000000000",  -- 27
	"000000000000000000000000",  -- 28
	"000000000000000000000000",  -- 29
	"000000000000000000000000",  -- 30
	"000000000000000000000000",  -- 31
--	"000000000000000000000000",  -- 32
--	"000011010000000000000000",  -- 32 -- JSR #0
	"000010111111000010000000",  -- 32 -- JSR absolute
	"000000000000000001000000",  -- 33 -- #64
	"000000000000000000000000",  -- 34
	"000000000000000000000000",  -- 35
	"000000000000000000000000",  -- 36
	"000000000000000000000000",  -- 37
	"000000000000000000000000",  -- 38
	"000000000000000000000000",  -- 39
	"000000000000000000000000",  -- 40
	"000000000000000000000000",  -- 41
	"000000000000000000000000",  -- 42
	"000000000000000000000000",  -- 43
	"000000000000000000000000",  -- 44
	"000000000000000000000000",  -- 45
	"000000000000000000000000",  -- 46
	"000000000000000000000000",  -- 47
	"000000000000000000000000",  -- 48
	"000000000000000000000000",  -- 49
	"000000000000000000000000",  -- 50
	"000000000000000000000000",  -- 51
	"000000000000000000000000",  -- 52
	"000000000000000000000000",  -- 53
	"000000000000000000000000",  -- 54
	"000000000000000000000000",  -- 55
	"000000000000000000000000",  -- 56
	"000000000000000000000000",  -- 57
	"000000000000000000000000",  -- 58
	"000000000000000000000000",  -- 59
	"000000000000000000000000",  -- 60
	"000000000000000000000000",  -- 61
	"000000000000000000000000",  -- 62
	"000000000000000000000000",  -- 63
	"000000000000000000000000",  -- 64
	"000000000000000000000000",  -- 65
	"000000000000000000000000",  -- 66
	"000000000000000000000000",  -- 67
	"000000000000000000000000",  -- 68
	"000000000000000000000000",  -- 69
	"000000000000000000000100",  -- 70 -- RTI
	"000000000000000000000000",  -- 71
	"000000000000000000000000",  -- 72
	"000000000000000000000000",  -- 73
	"000000000000000000000000",  -- 74
	"000000000000000000000000",  -- 75
	"000000000000000000000000",  -- 76
	"000000000000000000000000",  -- 77
	"000000000000000000000000",  -- 78
	"000000000000000000000000",  -- 79
	"000000000000000000000000",  -- 80
	"000000000000000000000000",  -- 81
	"000000000000000000000000",  -- 82
	"000000000000000000000000",  -- 83
	"000000000000000000000000",  -- 84
	"000000000000000000000000",  -- 85
	"000000000000000000000000",  -- 86
	"000000000000000000000000",  -- 87
	"000000000000000000000000",  -- 88
	"000000000000000000000000",  -- 89
	"000000000000000000000000",  -- 90
	"000000000000000000000000",  -- 91
	"000000000000000000000000",  -- 92
	"000000000000000000000000",  -- 93
	"000000000000000000000000",  -- 94
	"000000000000000000000000",  -- 95
	"000000000000000000000000",  -- 96
	"000000000000000000000000",  -- 97
	"000000000000000000000000",  -- 98
	"000000000000000000000000",  -- 99
	"000000000000000000000000",  -- 100
	"000000000000000000000000",  -- 101
	"000000000000000000000000",  -- 102
	"000000000000000000000000",  -- 103
	"000000000000000000000000",  -- 104
	"000000000000000000000000",  -- 105
	"000000000000000000000000",  -- 106
	"000000000000000000000000",  -- 107
	"000000000000000000000000",  -- 108
	"000000000000000000000000",  -- 109
	"000000000000000000000000",  -- 110
	"000000000000000000000000",  -- 111
	"000000000000000000000000",  -- 112
	"000000000000000000000000",  -- 113
	"000000000000000000000000",  -- 114
	"000000000000000000000000",  -- 115
	"000000000000000000000000",  -- 116
	"000000000000000000000000",  -- 117
	"000000000000000000000000",  -- 118
	"000000000000000000000000",  -- 119
	"000000000000000000000000",  -- 120
	"000000000000000000000000",  -- 121
	"000000000000000000000000",  -- 122
	"000000000000000000000000",  -- 123
	"000000000000000000000000",  -- 124
	"000000000000000000000000",  -- 125
	"000000000000000000000000",  -- 126
	"000000000000000000000000",  -- 127
	"000000000000000000000000",  -- 128
	"000000000000000000000000",  -- 129
	"000000000000000000000000",  -- 130
	"000000000000000000000000",  -- 131
	"000000000000000000000000",  -- 132
	"000000000000000000000000",  -- 133
	"000000000000000000000000",  -- 134
	"000000000000000000000000",  -- 135
	"000000000000000000000000",  -- 136
	"000000000000000000000000",  -- 137
	"000000000000000000000000",  -- 138
	"000000000000000000000000",  -- 139
	"000000000000000000000000",  -- 140
	"000000000000000000000000",  -- 141
	"000000000000000000000000",  -- 142
	"000000000000000000000000",  -- 143
	"000000000000000000000000",  -- 144
	"000000000000000000000000",  -- 145
	"000000000000000000000000",  -- 146
	"000000000000000000000000",  -- 147
	"000000000000000000000000",  -- 148
	"000000000000000000000000",  -- 149
	"000000000000000000000000",  -- 150
	"000000000000000000000000",  -- 151
	"000000000000000000000000",  -- 152
	"000000000000000000000000",  -- 153
	"000000000000000000000000",  -- 154
	"000000000000000000000000",  -- 155
	"000000000000000000000000",  -- 156
	"000000000000000000000000",  -- 157
	"000000000000000000000000",  -- 158
	"000000000000000000000000",  -- 159
	"000000000000000000000000",  -- 160
	"000000000000000000000000",  -- 161
	"000000000000000000000000",  -- 162
	"000000000000000000000000",  -- 163
	"000000000000000000000000",  -- 164
	"000000000000000000000000",  -- 165
	"000000000000000000000000",  -- 166
	"000000000000000000000000",  -- 167
	"000000000000000000000000",  -- 168
	"000000000000000000000000",  -- 169
	"000000000000000000000000",  -- 170
	"000000000000000000000000",  -- 171
	"000000000000000000000000",  -- 172
	"000000000000000000000000",  -- 173
	"000000000000000000000000",  -- 174
	"000000000000000000000000",  -- 175
	"000000000000000000000000",  -- 176
	"000000000000000000000000",  -- 177
	"000000000000000000000000",  -- 178
	"000000000000000000000000",  -- 179
	"000000000000000000000000",  -- 180
	"000000000000000000000000",  -- 181
	"000000000000000000000000",  -- 182
	"000000000000000000000000",  -- 183
	"000000000000000000000000",  -- 184
	"000000000000000000000000",  -- 185
	"000000000000000000000000",  -- 186
	"000000000000000000000000",  -- 187
	"000000000000000000000000",  -- 188
	"000000000000000000000000",  -- 189
	"000000000000000000000000",  -- 190
	"000000000000000000000000",  -- 191
	"000000000000000000000000",  -- 192
	"000000000000000000000000",  -- 193
	"000000000000000000000000",  -- 194
	"000000000000000000000000",  -- 195
	"000000000000000000000000",  -- 196
	"000000000000000000000000",  -- 197
	"000000000000000000000000",  -- 198
	"000000000000000000000000",  -- 199
	"000000000000000000000000",  -- 200
	"000000000000000000000000",  -- 201
	"000000000000000000000000",  -- 202
	"000000000000000000000000",  -- 203
	"000000000000000000000000",  -- 204
	"000000000000000000000000",  -- 205
	"000000000000000000000000",  -- 206
	"000000000000000000000000",  -- 207
	"000000000000000000000000",  -- 208
	"000000000000000000000000",  -- 209
	"000000000000000000000000",  -- 210
	"000000000000000000000000",  -- 211
	"000000000000000000000000",  -- 212
	"000000000000000000000000",  -- 213
	"000000000000000000000000",  -- 214
	"000000000000000000000000",  -- 215
	"000000000000000000000000",  -- 216
	"000000000000000000000000",  -- 217
	"000000000000000000000000",  -- 218
	"000000000000000000000000",  -- 219
	"000000000000000000000000",  -- 220
	"000000000000000000000000",  -- 221
	"000000000000000000000000",  -- 222
	"000000000000000000000000",  -- 223
	"000000000000000000000000",  -- 224
	"000000000000000000000000",  -- 225
	"000000000000000000000000",  -- 226
	"000000000000000000000000",  -- 227
	"000000000000000000000000",  -- 228
	"000000000000000000000000",  -- 229
	"000000000000000000000000",  -- 230
	"000000000000000000000000",  -- 231
	"000000000000000000000000",  -- 232
	"000000000000000000000000",  -- 233
	"000000000000000000000000",  -- 234
	"000000000000000000000000",  -- 235
	"000000000000000000000000",  -- 236
	"000000000000000000000000",  -- 237
	"000000000000000000000000",  -- 238
	"000000000000000000000000",  -- 239
	"000000000000000000000000",  -- 240
	"000000000000000000000000",  -- 241
	"000000000000000000000000",  -- 242
	"000000000000000000000000",  -- 243
	"000000000000000000000000",  -- 244
	"000000000000000000000000",  -- 245
	"000000000000000000000000",  -- 246
	"000000000000000000000000",  -- 247
	"000000000000000000000000",  -- 248
	"000000000000000000000000",  -- 249
	"000000000000000000000000",  -- 250
	"000000000000000000000000",  -- 251
	"000000000000000000000000",  -- 252
	"000000000000000000000000",  -- 253
	"000000000000000000000000",  -- 254
	"000000000000000000000000");  -- 255
	signal int_xmem : int_mem_type := (
--						when "11------10000000" => instr_array(JMP_INSTR)  <= '1';
--	"000000000000111011111001",  -- 0 -- ORI #$0E, CCR
	"000000000000000000001100",  -- 0 -- REP
	"000000000000000000000101",  -- 1 -- ORI #$0E, MR
	"000000000000111011111010",  -- 2 -- ORI #$0E, OMR
	"000000000000100010111010",  -- 3 -- ANDI #$08, OMR
--	"000010101111000010000000",  -- 1 -- JMP absolute
--	"000000000000000000011111",  -- 2 -- #31
--	"000011000000000000010000",  -- 3 -- JMP #16
	"000000000000000000000000",  -- 4
	"000000000000000000000000",  -- 5
	"000000000000000000000000",  -- 6
	"000000000000000000000000",  -- 7
	"000000000000000000000000",  -- 8
	"000000000000000000000000",  -- 9
	"000000000000000000000000",  -- 10
	"000000000000000000000000",  -- 11
	"000000000000000000000000",  -- 12
	"000000000000000000000000",  -- 13
	"000000000000000000000000",  -- 14
	"000000000000000000000000",  -- 15
	"000000000000000000000000",  -- 16
--	"000000000000000000000000",  -- 17
	"000010101101010110100000",  -- 17 -- JCC (r5)-
	"000000000000000000000000",  -- 18
	"000000000000000000000000",  -- 19
	"000010101101101010000000",  -- 20 -- JMP (r2)+
	"000000000000000000000000",  -- 21
	"000000000000000000000000",  -- 22
	"000000000000000000000000",  -- 23
	"000000000000000000000000",  -- 24
	"000000000000000000000000",  -- 25
	"000000000000000000000000",  -- 26
	"000000000000000000000000",  -- 27
	"000000000000000000000000",  -- 28
	"000000000000000000000000",  -- 29
	"000000000000000000000000",  -- 30
	"000000000000000000000000",  -- 31
--	"000000000000000000000000",  -- 32
--	"000011010000000000000000",  -- 32 -- JSR #0
	"000010111111000010000000",  -- 32 -- JSR absolute
	"000000000000000001000000",  -- 33 -- #64
	"000000000000000000000000",  -- 34
	"000000000000000000000000",  -- 35
	"000000000000000000000000",  -- 36
	"000000000000000000000000",  -- 37
	"000000000000000000000000",  -- 38
	"000000000000000000000000",  -- 39
	"000000000000000000000000",  -- 40
	"000000000000000000000000",  -- 41
	"000000000000000000000000",  -- 42
	"000000000000000000000000",  -- 43
	"000000000000000000000000",  -- 44
	"000000000000000000000000",  -- 45
	"000000000000000000000000",  -- 46
	"000000000000000000000000",  -- 47
	"000000000000000000000000",  -- 48
	"000000000000000000000000",  -- 49
	"000000000000000000000000",  -- 50
	"000000000000000000000000",  -- 51
	"000000000000000000000000",  -- 52
	"000000000000000000000000",  -- 53
	"000000000000000000000000",  -- 54
	"000000000000000000000000",  -- 55
	"000000000000000000000000",  -- 56
	"000000000000000000000000",  -- 57
	"000000000000000000000000",  -- 58
	"000000000000000000000000",  -- 59
	"000000000000000000000000",  -- 60
	"000000000000000000000000",  -- 61
	"000000000000000000000000",  -- 62
	"000000000000000000000000",  -- 63
	"000000000000000000000000",  -- 64
	"000000000000000000000000",  -- 65
	"000000000000000000000000",  -- 66
	"000000000000000000000000",  -- 67
	"000000000000000000000000",  -- 68
	"000000000000000000000000",  -- 69
	"000000000000000000000100",  -- 70 -- RTI
	"000000000000000000000000",  -- 71
	"000000000000000000000000",  -- 72
	"000000000000000000000000",  -- 73
	"000000000000000000000000",  -- 74
	"000000000000000000000000",  -- 75
	"000000000000000000000000",  -- 76
	"000000000000000000000000",  -- 77
	"000000000000000000000000",  -- 78
	"000000000000000000000000",  -- 79
	"000000000000000000000000",  -- 80
	"000000000000000000000000",  -- 81
	"000000000000000000000000",  -- 82
	"000000000000000000000000",  -- 83
	"000000000000000000000000",  -- 84
	"000000000000000000000000",  -- 85
	"000000000000000000000000",  -- 86
	"000000000000000000000000",  -- 87
	"000000000000000000000000",  -- 88
	"000000000000000000000000",  -- 89
	"000000000000000000000000",  -- 90
	"000000000000000000000000",  -- 91
	"000000000000000000000000",  -- 92
	"000000000000000000000000",  -- 93
	"000000000000000000000000",  -- 94
	"000000000000000000000000",  -- 95
	"000000000000000000000000",  -- 96
	"000000000000000000000000",  -- 97
	"000000000000000000000000",  -- 98
	"000000000000000000000000",  -- 99
	"000000000000000000000000",  -- 100
	"000000000000000000000000",  -- 101
	"000000000000000000000000",  -- 102
	"000000000000000000000000",  -- 103
	"000000000000000000000000",  -- 104
	"000000000000000000000000",  -- 105
	"000000000000000000000000",  -- 106
	"000000000000000000000000",  -- 107
	"000000000000000000000000",  -- 108
	"000000000000000000000000",  -- 109
	"000000000000000000000000",  -- 110
	"000000000000000000000000",  -- 111
	"000000000000000000000000",  -- 112
	"000000000000000000000000",  -- 113
	"000000000000000000000000",  -- 114
	"000000000000000000000000",  -- 115
	"000000000000000000000000",  -- 116
	"000000000000000000000000",  -- 117
	"000000000000000000000000",  -- 118
	"000000000000000000000000",  -- 119
	"000000000000000000000000",  -- 120
	"000000000000000000000000",  -- 121
	"000000000000000000000000",  -- 122
	"000000000000000000000000",  -- 123
	"000000000000000000000000",  -- 124
	"000000000000000000000000",  -- 125
	"000000000000000000000000",  -- 126
	"000000000000000000000000",  -- 127
	"000000000000000000000000",  -- 128
	"000000000000000000000000",  -- 129
	"000000000000000000000000",  -- 130
	"000000000000000000000000",  -- 131
	"000000000000000000000000",  -- 132
	"000000000000000000000000",  -- 133
	"000000000000000000000000",  -- 134
	"000000000000000000000000",  -- 135
	"000000000000000000000000",  -- 136
	"000000000000000000000000",  -- 137
	"000000000000000000000000",  -- 138
	"000000000000000000000000",  -- 139
	"000000000000000000000000",  -- 140
	"000000000000000000000000",  -- 141
	"000000000000000000000000",  -- 142
	"000000000000000000000000",  -- 143
	"000000000000000000000000",  -- 144
	"000000000000000000000000",  -- 145
	"000000000000000000000000",  -- 146
	"000000000000000000000000",  -- 147
	"000000000000000000000000",  -- 148
	"000000000000000000000000",  -- 149
	"000000000000000000000000",  -- 150
	"000000000000000000000000",  -- 151
	"000000000000000000000000",  -- 152
	"000000000000000000000000",  -- 153
	"000000000000000000000000",  -- 154
	"000000000000000000000000",  -- 155
	"000000000000000000000000",  -- 156
	"000000000000000000000000",  -- 157
	"000000000000000000000000",  -- 158
	"000000000000000000000000",  -- 159
	"000000000000000000000000",  -- 160
	"000000000000000000000000",  -- 161
	"000000000000000000000000",  -- 162
	"000000000000000000000000",  -- 163
	"000000000000000000000000",  -- 164
	"000000000000000000000000",  -- 165
	"000000000000000000000000",  -- 166
	"000000000000000000000000",  -- 167
	"000000000000000000000000",  -- 168
	"000000000000000000000000",  -- 169
	"000000000000000000000000",  -- 170
	"000000000000000000000000",  -- 171
	"000000000000000000000000",  -- 172
	"000000000000000000000000",  -- 173
	"000000000000000000000000",  -- 174
	"000000000000000000000000",  -- 175
	"000000000000000000000000",  -- 176
	"000000000000000000000000",  -- 177
	"000000000000000000000000",  -- 178
	"000000000000000000000000",  -- 179
	"000000000000000000000000",  -- 180
	"000000000000000000000000",  -- 181
	"000000000000000000000000",  -- 182
	"000000000000000000000000",  -- 183
	"000000000000000000000000",  -- 184
	"000000000000000000000000",  -- 185
	"000000000000000000000000",  -- 186
	"000000000000000000000000",  -- 187
	"000000000000000000000000",  -- 188
	"000000000000000000000000",  -- 189
	"000000000000000000000000",  -- 190
	"000000000000000000000000",  -- 191
	"000000000000000000000000",  -- 192
	"000000000000000000000000",  -- 193
	"000000000000000000000000",  -- 194
	"000000000000000000000000",  -- 195
	"000000000000000000000000",  -- 196
	"000000000000000000000000",  -- 197
	"000000000000000000000000",  -- 198
	"000000000000000000000000",  -- 199
	"000000000000000000000000",  -- 200
	"000000000000000000000000",  -- 201
	"000000000000000000000000",  -- 202
	"000000000000000000000000",  -- 203
	"000000000000000000000000",  -- 204
	"000000000000000000000000",  -- 205
	"000000000000000000000000",  -- 206
	"000000000000000000000000",  -- 207
	"000000000000000000000000",  -- 208
	"000000000000000000000000",  -- 209
	"000000000000000000000000",  -- 210
	"000000000000000000000000",  -- 211
	"000000000000000000000000",  -- 212
	"000000000000000000000000",  -- 213
	"000000000000000000000000",  -- 214
	"000000000000000000000000",  -- 215
	"000000000000000000000000",  -- 216
	"000000000000000000000000",  -- 217
	"000000000000000000000000",  -- 218
	"000000000000000000000000",  -- 219
	"000000000000000000000000",  -- 220
	"000000000000000000000000",  -- 221
	"000000000000000000000000",  -- 222
	"000000000000000000000000",  -- 223
	"000000000000000000000000",  -- 224
	"000000000000000000000000",  -- 225
	"000000000000000000000000",  -- 226
	"000000000000000000000000",  -- 227
	"000000000000000000000000",  -- 228
	"000000000000000000000000",  -- 229
	"000000000000000000000000",  -- 230
	"000000000000000000000000",  -- 231
	"000000000000000000000000",  -- 232
	"000000000000000000000000",  -- 233
	"000000000000000000000000",  -- 234
	"000000000000000000000000",  -- 235
	"000000000000000000000000",  -- 236
	"000000000000000000000000",  -- 237
	"000000000000000000000000",  -- 238
	"000000000000000000000000",  -- 239
	"000000000000000000000000",  -- 240
	"000000000000000000000000",  -- 241
	"000000000000000000000000",  -- 242
	"000000000000000000000000",  -- 243
	"000000000000000000000000",  -- 244
	"000000000000000000000000",  -- 245
	"000000000000000000000000",  -- 246
	"000000000000000000000000",  -- 247
	"000000000000000000000000",  -- 248
	"000000000000000000000000",  -- 249
	"000000000000000000000000",  -- 250
	"000000000000000000000000",  -- 251
	"000000000000000000000000",  -- 252
	"000000000000000000000000",  -- 253
	"000000000000000000000000",  -- 254
	"000000000000000000000000");  -- 255
	signal int_ymem : int_mem_type := (
--						when "11------10000000" => instr_array(JMP_INSTR)  <= '1';
--	"000000000000111011111001",  -- 0 -- ORI #$0E, CCR
	"000000000000000000000001",  -- 0 -- REP
	"000000000000000000000010",  -- 1 -- ORI #$0E, MR
	"000000000000000000000011",  -- 2 -- ORI #$0E, OMR
	"000000000000000000000100",  -- 3 -- ANDI #$08, OMR
--	"000010101111000010000000",  -- 1 -- JMP absolute
--	"000000000000000000011111",  -- 2 -- #31
--	"000011000000000000010000",  -- 3 -- JMP #16
	"000000000000000000000101",  -- 4
	"000000000000000000000110",  -- 5
	"000000000000000000000111",  -- 6
	"000000000000000000001000",  -- 7
	"000000000000000000001001",  -- 8
	"000000000000000000001010",  -- 9
	"000000000000000000001011",  -- 10
	"000000000000000000001100",  -- 11
	"000000000000000000001101",  -- 12
	"000000000000000000001110",  -- 13
	"000000000000000000001111",  -- 14
	"000000000000000000010000",  -- 15
	"000000000000000000010001",  -- 16
--	"000000000000000000000000",  -- 17
	"000010101101010110100000",  -- 17 -- JCC (r5)-
	"000000000000000000000000",  -- 18
	"000000000000000000000000",  -- 19
	"000010101101101010000000",  -- 20 -- JMP (r2)+
	"000000000000000000000000",  -- 21
	"000000000000000000000000",  -- 22
	"000000000000000000000000",  -- 23
	"000000000000000000000000",  -- 24
	"000000000000000000000000",  -- 25
	"000000000000000000000000",  -- 26
	"000000000000000000000000",  -- 27
	"000000000000000000000000",  -- 28
	"000000000000000000000000",  -- 29
	"000000000000000000000000",  -- 30
	"000000000000000000000000",  -- 31
--	"000000000000000000000000",  -- 32
--	"000011010000000000000000",  -- 32 -- JSR #0
	"000010111111000010000000",  -- 32 -- JSR absolute
	"000000000000000001000000",  -- 33 -- #64
	"000000000000000000000000",  -- 34
	"000000000000000000000000",  -- 35
	"000000000000000000000000",  -- 36
	"000000000000000000000000",  -- 37
	"000000000000000000000000",  -- 38
	"000000000000000000000000",  -- 39
	"000000000000000000000000",  -- 40
	"000000000000000000000000",  -- 41
	"000000000000000000000000",  -- 42
	"000000000000000000000000",  -- 43
	"000000000000000000000000",  -- 44
	"000000000000000000000000",  -- 45
	"000000000000000000000000",  -- 46
	"000000000000000000000000",  -- 47
	"000000000000000000000000",  -- 48
	"000000000000000000000000",  -- 49
	"000000000000000000000000",  -- 50
	"000000000000000000000000",  -- 51
	"000000000000000000000000",  -- 52
	"000000000000000000000000",  -- 53
	"000000000000000000000000",  -- 54
	"000000000000000000000000",  -- 55
	"000000000000000000000000",  -- 56
	"000000000000000000000000",  -- 57
	"000000000000000000000000",  -- 58
	"000000000000000000000000",  -- 59
	"000000000000000000000000",  -- 60
	"000000000000000000000000",  -- 61
	"000000000000000000000000",  -- 62
	"000000000000000000000000",  -- 63
	"000000000000000000000000",  -- 64
	"000000000000000000000000",  -- 65
	"000000000000000000000000",  -- 66
	"000000000000000000000000",  -- 67
	"000000000000000000000000",  -- 68
	"000000000000000000000000",  -- 69
	"000000000000000000000100",  -- 70 -- RTI
	"000000000000000000000000",  -- 71
	"000000000000000000000000",  -- 72
	"000000000000000000000000",  -- 73
	"000000000000000000000000",  -- 74
	"000000000000000000000000",  -- 75
	"000000000000000000000000",  -- 76
	"000000000000000000000000",  -- 77
	"000000000000000000000000",  -- 78
	"000000000000000000000000",  -- 79
	"000000000000000000000000",  -- 80
	"000000000000000000000000",  -- 81
	"000000000000000000000000",  -- 82
	"000000000000000000000000",  -- 83
	"000000000000000000000000",  -- 84
	"000000000000000000000000",  -- 85
	"000000000000000000000000",  -- 86
	"000000000000000000000000",  -- 87
	"000000000000000000000000",  -- 88
	"000000000000000000000000",  -- 89
	"000000000000000000000000",  -- 90
	"000000000000000000000000",  -- 91
	"000000000000000000000000",  -- 92
	"000000000000000000000000",  -- 93
	"000000000000000000000000",  -- 94
	"000000000000000000000000",  -- 95
	"000000000000000000000000",  -- 96
	"000000000000000000000000",  -- 97
	"000000000000000000000000",  -- 98
	"000000000000000000000000",  -- 99
	"000000000000000000000000",  -- 100
	"000000000000000000000000",  -- 101
	"000000000000000000000000",  -- 102
	"000000000000000000000000",  -- 103
	"000000000000000000000000",  -- 104
	"000000000000000000000000",  -- 105
	"000000000000000000000000",  -- 106
	"000000000000000000000000",  -- 107
	"000000000000000000000000",  -- 108
	"000000000000000000000000",  -- 109
	"000000000000000000000000",  -- 110
	"000000000000000000000000",  -- 111
	"000000000000000000000000",  -- 112
	"000000000000000000000000",  -- 113
	"000000000000000000000000",  -- 114
	"000000000000000000000000",  -- 115
	"000000000000000000000000",  -- 116
	"000000000000000000000000",  -- 117
	"000000000000000000000000",  -- 118
	"000000000000000000000000",  -- 119
	"000000000000000000000000",  -- 120
	"000000000000000000000000",  -- 121
	"000000000000000000000000",  -- 122
	"000000000000000000000000",  -- 123
	"000000000000000000000000",  -- 124
	"000000000000000000000000",  -- 125
	"000000000000000000000000",  -- 126
	"000000000000000000000000",  -- 127
	"000000000000000000000000",  -- 128
	"000000000000000000000000",  -- 129
	"000000000000000000000000",  -- 130
	"000000000000000000000000",  -- 131
	"000000000000000000000000",  -- 132
	"000000000000000000000000",  -- 133
	"000000000000000000000000",  -- 134
	"000000000000000000000000",  -- 135
	"000000000000000000000000",  -- 136
	"000000000000000000000000",  -- 137
	"000000000000000000000000",  -- 138
	"000000000000000000000000",  -- 139
	"000000000000000000000000",  -- 140
	"000000000000000000000000",  -- 141
	"000000000000000000000000",  -- 142
	"000000000000000000000000",  -- 143
	"000000000000000000000000",  -- 144
	"000000000000000000000000",  -- 145
	"000000000000000000000000",  -- 146
	"000000000000000000000000",  -- 147
	"000000000000000000000000",  -- 148
	"000000000000000000000000",  -- 149
	"000000000000000000000000",  -- 150
	"000000000000000000000000",  -- 151
	"000000000000000000000000",  -- 152
	"000000000000000000000000",  -- 153
	"000000000000000000000000",  -- 154
	"000000000000000000000000",  -- 155
	"000000000000000000000000",  -- 156
	"000000000000000000000000",  -- 157
	"000000000000000000000000",  -- 158
	"000000000000000000000000",  -- 159
	"000000000000000000000000",  -- 160
	"000000000000000000000000",  -- 161
	"000000000000000000000000",  -- 162
	"000000000000000000000000",  -- 163
	"000000000000000000000000",  -- 164
	"000000000000000000000000",  -- 165
	"000000000000000000000000",  -- 166
	"000000000000000000000000",  -- 167
	"000000000000000000000000",  -- 168
	"000000000000000000000000",  -- 169
	"000000000000000000000000",  -- 170
	"000000000000000000000000",  -- 171
	"000000000000000000000000",  -- 172
	"000000000000000000000000",  -- 173
	"000000000000000000000000",  -- 174
	"000000000000000000000000",  -- 175
	"000000000000000000000000",  -- 176
	"000000000000000000000000",  -- 177
	"000000000000000000000000",  -- 178
	"000000000000000000000000",  -- 179
	"000000000000000000000000",  -- 180
	"000000000000000000000000",  -- 181
	"000000000000000000000000",  -- 182
	"000000000000000000000000",  -- 183
	"000000000000000000000000",  -- 184
	"000000000000000000000000",  -- 185
	"000000000000000000000000",  -- 186
	"000000000000000000000000",  -- 187
	"000000000000000000000000",  -- 188
	"000000000000000000000000",  -- 189
	"000000000000000000000000",  -- 190
	"000000000000000000000000",  -- 191
	"000000000000000000000000",  -- 192
	"000000000000000000000000",  -- 193
	"000000000000000000000000",  -- 194
	"000000000000000000000000",  -- 195
	"000000000000000000000000",  -- 196
	"000000000000000000000000",  -- 197
	"000000000000000000000000",  -- 198
	"000000000000000000000000",  -- 199
	"000000000000000000000000",  -- 200
	"000000000000000000000000",  -- 201
	"000000000000000000000000",  -- 202
	"000000000000000000000000",  -- 203
	"000000000000000000000000",  -- 204
	"000000000000000000000000",  -- 205
	"000000000000000000000000",  -- 206
	"000000000000000000000000",  -- 207
	"000000000000000000000000",  -- 208
	"000000000000000000000000",  -- 209
	"000000000000000000000000",  -- 210
	"000000000000000000000000",  -- 211
	"000000000000000000000000",  -- 212
	"000000000000000000000000",  -- 213
	"000000000000000000000000",  -- 214
	"000000000000000000000000",  -- 215
	"000000000000000000000000",  -- 216
	"000000000000000000000000",  -- 217
	"000000000000000000000000",  -- 218
	"000000000000000000000000",  -- 219
	"000000000000000000000000",  -- 220
	"000000000000000000000000",  -- 221
	"000000000000000000000000",  -- 222
	"000000000000000000000000",  -- 223
	"000000000000000000000000",  -- 224
	"000000000000000000000000",  -- 225
	"000000000000000000000000",  -- 226
	"000000000000000000000000",  -- 227
	"000000000000000000000000",  -- 228
	"000000000000000000000000",  -- 229
	"000000000000000000000000",  -- 230
	"000000000000000000000000",  -- 231
	"000000000000000000000000",  -- 232
	"000000000000000000000000",  -- 233
	"000000000000000000000000",  -- 234
	"000000000000000000000000",  -- 235
	"000000000000000000000000",  -- 236
	"000000000000000000000000",  -- 237
	"000000000000000000000000",  -- 238
	"000000000000000000000000",  -- 239
	"000000000000000000000000",  -- 240
	"000000000000000000000000",  -- 241
	"000000000000000000000000",  -- 242
	"000000000000000000000000",  -- 243
	"000000000000000000000000",  -- 244
	"000000000000000000000000",  -- 245
	"000000000000000000000000",  -- 246
	"000000000000000000000000",  -- 247
	"000000000000000000000000",  -- 248
	"000000000000000000000000",  -- 249
	"000000000000000000000000",  -- 250
	"000000000000000000000000",  -- 251
	"000000000000000000000000",  -- 252
	"000000000000000000000000",  -- 253
	"000000000000000000000000",  -- 254
	"000000000000000000000000");  -- 255

begin

--	int_mem <= int_pmem when mem_type = P_MEM else
--	           int_xmem when mem_type = X_MEM else
--	           int_ymem when mem_type = Y_MEM;

	wr_accomplished <= wr_en;

	PMEM_GEN: if mem_type = P_MEM generate
		data_out <= int_pmem(to_integer(unsigned(int_mem_rd_addr)));
		process(clk) is
		begin
			if rising_edge(clk) then
--				if rst = '1' then
--					data_out_valid <= '0';
--					int_mem_rd_addr <= (others => '0');
--				else
					int_mem_rd_addr <= std_logic_vector(rd_addr(7 downto 0));
					data_out_valid <= rd_en;
					if wr_en = '1' then
							int_pmem(to_integer(wr_addr)) <= data_in;
					end if;
--				end if;
			end if;
		end process;
	end generate;

	XMEM_GEN: if mem_type = X_MEM generate
		data_out <= int_xmem(to_integer(unsigned(int_mem_rd_addr)));
		process(clk) is
		begin
			if rising_edge(clk) then
--				if rst = '1' then
--					data_out_valid <= '0';
--					int_mem_rd_addr <= (others => '0');
--				else
					int_mem_rd_addr <= std_logic_vector(rd_addr(7 downto 0));
					data_out_valid <= rd_en;
					if wr_en = '1' then
							int_xmem(to_integer(wr_addr)) <= data_in;
					end if;
--				end if;
			end if;
		end process;
	end generate;

	YMEM_GEN: if mem_type = Y_MEM generate
		data_out <= int_ymem(to_integer(unsigned(int_mem_rd_addr)));
		process(clk) is
		begin
			if rising_edge(clk) then
--				if rst = '1' then
--					data_out_valid <= '0';
--					int_mem_rd_addr <= (others => '0');
--				else
					int_mem_rd_addr <= std_logic_vector(rd_addr(7 downto 0));
					data_out_valid <= rd_en;
					if wr_en = '1' then
							int_ymem(to_integer(wr_addr)) <= data_in;
					end if;
--				end if;
			end if;
		end process;
	end generate;
--	process(clk, rst) is
--	begin
--		if rising_edge(clk) then
--			if rst = '1' then
--				data_out_valid <= '0';
--				int_mem_rd_addr <= (others => '0');
--			else
--				int_mem_rd_addr <= std_logic_vector(rd_addr(7 downto 0));
--				data_out_valid <= rd_en;
--				if wr_en = '1' then
--					if mem_type = P_MEM then
--						int_pmem(to_integer(wr_addr)) <= data_in;
--					elsif mem_type = X_MEM then
--						int_xmem(to_integer(wr_addr)) <= data_in;
--					elsif mem_type = Y_MEM then
--						int_ymem(to_integer(wr_addr)) <= data_in;
--					end if;
--				end if;
--			end if;
--		end if;
--	end process;

end architecture rtl;

