
package parameter_pkg is

	constant BW_ADDRESS : natural := 16;

	constant PIPELINE_DEPTH : natural := 5;

	constant NUM_ACT_SIGNALS : natural := 26;

end package;
